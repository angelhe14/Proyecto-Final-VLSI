library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity proyecto is

end proyecto;

architecture behavioral of proyecto is



end behavioral;